module Paraller_Multiplier (
	input logic [31:0] Multiplier,
	input logic [31:0] Multiplicand 
);


endmodule