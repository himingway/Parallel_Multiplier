module CompressTree (
	input logic [15:0] Error_Correction,
	input logic [33:0] PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, 
		PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15,
	input logic [31:0] PP16,
	output logic [63:0] C,
	output logic [63:0] S
);

logic ZERO;

assign ZERO = 0;

logic [33:0] C11; logic [33:0] S11; logic [33:0] C12; logic [33:0] S12;
logic [33:0] C13; logic [33:0] S13; logic [33:0] C14; logic [33:0] S14;
logic [33:0] C21; logic [33:0] S21; logic [37:0] C22; logic [37:0] S22;
logic [33:0] C23; logic [33:0] S23; logic [33:0] C24; logic [33:0] S24;
logic [39:0] C31; logic [39:0] S31; logic [38:0] C32; logic[38:0] S32;
logic [45:0] C41; logic [45:0] S41; logic [45:0] C42; logic[45:0] S42;
logic [46:0] C51; logic [46:0] S51; logic [56:0] C61; logic[56:0] S61;
logic [63:0] C71; logic [63:0] S71;

assign C = C71;
assign S = S71;

Carry_Save_Adder #34 CSA13(
	.a({{4{PP0[33]}}, PP0[33:4]}), 
	.b({{2{PP1[33]}}, PP1[33:2]}), 
	.Cin(PP2[33:0]), 
	.Cout(C13), .Sum(S13));

Carry_Save_Adder #34 CSA23(
	.a(PP3[33:0]), 
	.b({C13[33], C13[33:1]}), 
	.Cin({{2{S13[33]}}, S13[33:2]}), 
	.Cout(C23), .Sum(S23));

Carry_Save_Adder #34 CSA14(
	.a({{4{PP4[33]}}, PP4[33:4]}), 
	.b({{2{PP5[33]}}, PP5[33:2]}), 
	.Cin(PP6[33:0]), 
	.Cout(C14), .Sum(S14));

Carry_Save_Adder #34 CSA24(
	.a({{2{PP7[33]}}, PP7[33:2]}), 
	.b(PP8[33:0]), 
	.Cin({{3{C14[33]}}, C14[33:3]}), 
	.Cout(C24), .Sum(S24));

Carry_Save_Adder #34 CSA11(
	.a({{4{PP9[33]}}, PP9[33:4]}), 
	.b({{2{PP10[33]}}, PP10[33:2]}), 
	.Cin(PP11[33:0]), 
	.Cout(C11), .Sum(S11));

Carry_Save_Adder #34 CSA21(
	.a(PP12[33:0]), 
	.b({C11[33], C11[33:1]}), 
	.Cin({{2{S11[33]}}, S11[33:2]}), 
	.Cout(C21), .Sum(S21));

Carry_Save_Adder #34 CSA12(
	.a({{4{PP13[33]}}, PP13[33:4]}), 
	.b({{2{PP14[33]}}, PP14[33:2]}), 
	.Cin(PP15[33:0]), 
	.Cout(C12), .Sum(S12));

Carry_Save_Adder #38 CSA22(
	.a({PP16[31:0], ZERO, Error_Correction[15], {PP13[3:0]}}), 
	.b({C12[32:0], ZERO, {PP14[1:0], {2{ZERO}}}}), 
	.Cin({S12[33:0], ZERO, Error_Correction[14], ZERO, Error_Correction[13]}), 
	.Cout(C22), .Sum(S22));

Carry_Save_Adder #40 CSA31(
	.a({{6{S21[33]}}, S21[33:0]}), 
	.b({C22[36:0], {3{ZERO}}}), 
	.Cin({S22[37:0], ZERO, Error_Correction[12]}), 
	.Cout(C31), .Sum(S31));

Carry_Save_Adder #39 CSA32(
	.a({C24[33:0], ZERO, {PP7[1:0], ZERO}, ZERO}), 
	.b({S24[33], S24[33:0], {C14[2:0]}, ZERO}), 
	.Cin({{5{S14[33]}}, S14[33:0]}), 
	.Cout(C32), .Sum(S32));

Carry_Save_Adder #46 CSA41(
	.a({{5{C21[33]}}, C21[33:0], ZERO, {C11[0], ZERO}, {PP9[3:0]}}), 
	.b({C31[38:0], ZERO, {S11[1:0]}, {PP10[1:0], {2{ZERO}}}}), 
	.Cin({S31[39:0], ZERO, Error_Correction[11], ZERO, Error_Correction[10], ZERO, Error_Correction[9]}), 
	.Cout(C41), .Sum(S41));

Carry_Save_Adder #46 CSA42(
	.a({{11{C23[33]}}, C23[33:0], ZERO}), 
	.b({{12{S23[33]}}, S23[33:0]}), 
	.Cin({C32[38:0], Error_Correction[6], ZERO, Error_Correction[5], ZERO, Error_Correction[4], ZERO, Error_Correction[3]}), 
	.Cout(C42), .Sum(S42));

Carry_Save_Adder #47 CSA51(
	.a({C42[45:0], ZERO}), 
	.b({{2{S32[38]}}, S32[38:0], {6{ZERO}}}), 
	.Cin({S42[45], S42[45:0]}), 
	.Cout(C51), .Sum(S51));

Carry_Save_Adder #57 CSA61(
	.a({C41[44:0], {7{ZERO}}, {PP4[3:0]}, ZERO}), 
	.b({S41[45:0], ZERO, Error_Correction[8], ZERO, Error_Correction[7], {2{ZERO}}, {PP5[1:0], {2{ZERO}}}, ZERO}), 
	.Cin({{10{C51[46]}}, C51[46:0]}), 
	.Cout(C61), .Sum(S61));

Carry_Save_Adder #64 CSA71(
	.a({C61[55:0], {2{ZERO}}, {C13[0], ZERO}, {PP0[3:0]}}), 
	.b({S61[56:0], ZERO, {S13[1:0]}, {PP1[1:0], {2{ZERO}}}}), 
	.Cin({{11{S51[46]}}, S51[46:0], ZERO, Error_Correction[2], ZERO, Error_Correction[1], ZERO, Error_Correction[0]}), 
	.Cout(C71), .Sum(S71));

endmodule